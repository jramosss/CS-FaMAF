/*
Realizar un testbench usando señales de entrada que permitan, a partir del análisis de las salidas
resultantes, verificar la correcta instanciación y conexionado de todos los módulos y caminos de
señal de la estructura interna del módulo execute.
*/
module execute_tb ();
	
endmodule 