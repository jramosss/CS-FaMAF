//- Ingrese por el puerto a todos los tipos de instrucciones detalladas en la tabla, con
//inmediatos positivos y negativos, y verifique que la salida sea la correcta.
//- Ingrese instrucciones que no estén en la tabla y verifique que la salida sea 0

/*
module signext_tb();
	logic lit = 0;
	logic LDUR = 
	
*/